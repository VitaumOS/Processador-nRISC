library verilog;
use verilog.vl_types.all;
entity nRisc_Simula is
end nRisc_Simula;
