module Somador(
	
	input wire [7:0] d1,d2,
	
	output reg [7:0] saida
);

	always @* begin
	
		saida = d1+d2;
	end

endmodule
